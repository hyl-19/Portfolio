module DFF(q, d, clk, reset);

  output q; 
  input d, clk, reset;
  reg q;

  always @(posedge reset or negedge clk) 
    if (reset)
		    q = 1'b0;
    else
		    q = d;


endmodule
//========================================
module MUX4_1(s0, s1, i0, i1, i2, i3, out);
  output out ;
  input s0, s1, i0, i1, i2, i3;
  
  assign out = s1 ? ( s0 ? i3 : i2 ) :( s0 ? i1 : i0 ) ;
  
endmodule
//========================================
module Shift_Register(i ,s ,o ,clk, reset, r);
  output[7:0] o; 
  input[7:0] i;
  input[1:0] s;
  input r, clk, reset;
  reg[7:0] o;
  wire a0, a1, a2, a3, a4, a5, a6, a7 ;
  wire mo0, mo1, mo2, mo3, mo4, mo5, mo6, mo7; // out of mux
  
    MUX4_1 M0( s[0], s[1], a0, r , a1, i[0], mo0 );
    MUX4_1 M1( s[0], s[1], a1, a0, a2, i[1], mo1 );
    MUX4_1 M2( s[0], s[1], a2, a1, a3, i[2], mo2 );
    MUX4_1 M3( s[0], s[1], a3, a2, a4, i[3], mo3 );
    MUX4_1 M4( s[0], s[1], a4, a3, a5, i[4], mo4 );
    MUX4_1 M5( s[0], s[1], a5, a4, a6, i[5], mo5 );
    MUX4_1 M6( s[0], s[1], a6, a5, a7, i[6], mo6 );
    MUX4_1 M7( s[0], s[1], a7, a6, r , i[7], mo7 );
    
    DFF D0(a0, mo0, clk, reset);
    DFF D1(a1, mo1, clk, reset);
    DFF D2(a2, mo2, clk, reset);
    DFF D3(a3, mo3, clk, reset);
    DFF D4(a4, mo4, clk, reset);
    DFF D5(a5, mo5, clk, reset);
    DFF D6(a6, mo6, clk, reset);
    DFF D7(a7, mo7, clk, reset);
    
  always @(posedge reset or negedge clk)
  if(reset)
    assign o = 8'b0000000;
  else 
    assign o = {a7, a6, a5, a4, a3, a2, a1, a0} ;
    
endmodule







