library verilog;
use verilog.vl_types.all;
entity tb_pipelined is
end tb_pipelined;
